#CUI|TUI|CODE|SAB|STR|PREF
C0027424|T184|68235000|SNOMEDCT_US|Nasal congestion|Congestion or runny nose
C1260880|T184|64531003|SNOMEDCT_US|Rhinorrhea|Congestion or runny nose
C0010200|T184|49727002|SNOMEDCT_US|Coughing|Cough
C0850149|T184|11833005|SNOMEDCT_US|Dry Cough|Cough
C0239134|T033|28743005|SNOMEDCT_US|Productive Cough|Cough
C0011991|T184|62315008|SNOMEDCT_US|Diarrhea|Diarrhea
C0015672|T184|84229001|SNOMEDCT_US|Fatigue|Fatigue
C0231218|T184|367391008|SNOMEDCT_US|Malaise|Fatigue
C0085593|T184|43724002|SNOMEDCT_US|Chills|Fever or chills
C0036973|T033|43724002|SNOMEDCT_US|Shivering|Fever or chills
C0687681|T184|103001002|SNOMEDCT_US|Feeling feverish|Fever or chills
C1959900|T033|426000000|SNOMEDCT_US|Fever greater than 100.4 Fahrenheit|Fever or chills
C0015967|T184|386661006|SNOMEDCT_US|Fever|Fever or chills
C0085594|T184|274640006|SNOMEDCT_US|Fever with chills|Fever or chills
C0018681|T184|25064002|SNOMEDCT_US|Headache|Headache
C0231528|T184|68962001|SNOMEDCT_US|Myalgia|Muscle or body aches
C0281856|T184|82991003|SNOMEDCT_US|Generalized aches and pains|Muscle or body aches
C0027497|T184|422587007|SNOMEDCT_US|Nausea|Nausea or vomiting
C0042963|T184|422400008|SNOMEDCT_US|Vomiting|Nausea or vomiting
C0027498|T184|16932000|SNOMEDCT_US|Nausea and vomiting|Nausea or vomiting
C0003126|T033|44169009|SNOMEDCT_US|Anosmia|Anosmia
C2364111|T184|36955009|SNOMEDCT_US|Ageusia|Anosmia
C0013378|T033|36955009|SNOMEDCT_US|Dysgeusia|Anosmia
C0013404|T184|267036007|SNOMEDCT_US|Dyspnea|Dyspnea
C0242429|T184|162397003|SNOMEDCT_US|Sore throat|Sore throat