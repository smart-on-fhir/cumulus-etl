#CUI|CODE|SAB|STR|PREF
C0027424|68235000|SNOMEDCT_US|Nasal congestion|Congestion or runny nose
C1260880|64531003|SNOMEDCT_US|Rhinorrhea|Congestion or runny nose
C0010200|49727002|SNOMEDCT_US|Coughing|Cough
C0850149|11833005|SNOMEDCT_US|Dry Cough|Cough
C0239134|28743005|SNOMEDCT_US|Productive Cough|Cough
C0011991|62315008|SNOMEDCT_US|Diarrhea|Diarrhea
C0015672|84229001|SNOMEDCT_US|Fatigue|Fatigue
C0231218|367391008|SNOMEDCT_US|Malaise|Fatigue
C0085593|43724002|SNOMEDCT_US|Chills|Fever or chills
C0036973|43724002|SNOMEDCT_US|Shivering|Fever or chills
C0687681|103001002|SNOMEDCT_US|Feeling feverish|Fever or chills
C1959900|426000000|SNOMEDCT_US|Fever greater than 100.4 Fahrenheit|Fever or chills
C0015967|386661006|SNOMEDCT_US|Fever|Fever or chills
C0085594|274640006|SNOMEDCT_US|Fever with chills|Fever or chills
C0018681|25064002|SNOMEDCT_US|Headache|Headache
C0231528|68962001|SNOMEDCT_US|Myalgia|Muscle or body aches
C0281856|82991003|SNOMEDCT_US|Generalized aches and pains|Muscle or body aches
C0027497|422587007|SNOMEDCT_US|Nausea|Nausea or vomiting
C0042963|422400008|SNOMEDCT_US|Vomiting|Nausea or vomiting
C0027498|16932000|SNOMEDCT_US|Nausea and vomiting|Nausea or vomiting
C0003126|44169009|SNOMEDCT_US|Anosmia|Anosmia
C2364111|36955009|SNOMEDCT_US|Ageusia|Anosmia
C0013378|36955009|SNOMEDCT_US|Dysgeusia|Anosmia
C0013404|267036007|SNOMEDCT_US|Dyspnea|Shortness of breath or difficulty breathing
C0242429|162397003|SNOMEDCT_US|Sore throat|Sore throat